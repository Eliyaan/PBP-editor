module pbp_g2c

// graph to code

const letters = ['a', 'b', 'c', 'd', 'e', 'f', 'g', 'h', 'i', 'j', 'k', 'l', 'm', 'n', 'o', 'p']

pub interface Graph {
	// blocks
	b_inps [][]int  // index of the ports
	b_outs [][]int  // index of the ports
	b_name []string // name of the block // fn names
	// ports
	p_input []bool   // is input or output
	p_name  []string // type names
	p_block []int    // index of block
	p_link  [][]int  // index of link
	// links
	l_inp []int // index of the input port
	l_out []int
}

pub fn generate_code(g Graph) string {
	mut output := '// AUTOGENERATED by pbp_editor\n'

	// import
	output += 'import pbp\n'
	output += 'import sync.stdatomic as atom\n'
	output += 'import runtime\n'

	// main
	// init queues (one for each input)
	output += 'fn main() {\n'
	for i, is_input in g.p_input {
		if is_input {
			output += '\tmut inp_${i}_${g.b_name[g.p_block[i]]} := pbp.AtomicQueue[${g.p_name[i]}]{}\n'
		}
	}
	output += '\tmut parts := []pbp.Part{}\n'
	// init the parts (one for each block)
	for i, name in g.b_name {
		name_camel_case := name.snake_to_camel()
		output += '\tparts << ${name_camel_case}{\n'
		for j, inp in g.b_inps[i] {
			output += '\t\t${letters[j]}_in: &inp_${inp}_${name}\n'
		}
		for j, out in g.b_outs[i] {
			output += '\t\t${letters[j]}_out: pbp.FanOut[${g.p_name[out]}]{['
			// links
			for k, link in g.p_link[out] {
				output += '&inp_${g.l_out[link]}_${g.b_name[g.p_block[g.l_out[link]]]}'
				if k != g.p_link[out].len - 1 {
					output += ', '
				}
			}
			output += ']}\n'
		}
		output += '\t}\n'
	}
	output += '\n\n'

	// run the threads
	output += '\tmut ths := []thread{}\n'
	output += '\tfor _ in 0 .. runtime.nr_cpus() {\n'
	output += '\t\tths << spawn pbp.part_runner(mut parts)\n'
	output += '\t}\n'
	output += '\tths.wait()\n'

	output += '}\n\n'

	for i, name in g.b_name {
		// fn struct
		name_camel_case := name.snake_to_camel()
		output += 'struct ' + name_camel_case + ' {\n'
		output += '\tf fn ('
		for j, inp in g.b_inps[i] {
			output += letters[j] + ' ' + g.p_name[inp]
			if j != g.b_inps[i].len - 1 {
				output += ','
			}
		}
		output += ') '
		if g.b_outs.len > 1 {
			output += '('
		}
		for j, out in g.b_outs[i] {
			output += ' ' + g.p_name[out]
			if j != g.b_outs[i].len - 1 {
				output += ','
			}
		}
		if g.b_outs.len > 1 {
			output += ')'
		}
		output += ' = ' + name + '\n'

		output += 'mut:\n'
		output += '\tready &atom.AtomicVal[bool] = atom.new_atomic(true)\n'

		for j, inp in g.b_inps[i] {
			output += '\t${letters[j]}_in &pbp.AtomicQueue[${inp}]\n'
		}
		for j, out in g.b_outs[i] {
			output += '\t${letters[j]}_out pbp.FanOut[${out}]\n'
		}
		output += '}\n\n'

		// run fn	
		output += 'fn (mut a ${name_camel_case}) run() {\n'
		output += '\tif '
		for j, _ in g.b_inps[i] {
			output += '!a.${letters[j]}_in.is_empty() '
			if j != g.b_inps[i].len - 1 {
				output += '&& '
			}
		}
		output += '{\n'
		// pop all the inputs from the queues
		for j, _ in g.b_inps[i] {
			l := letters[j]
			output += '\t\t${l}_in := a.${l}_in.pop() or { panic(@LOCATION) }\n'
		}
		// get all the outputs
		output += '\t\t'
		for j, _ in g.b_outs[i] {
			l := letters[j]
			output += l + '_out'
			if j != g.b_outs[i].len - 1 {
				output += ', '
			}
		}
		if g.b_outs[i].len >= 1 {
			output += ' := '
		}
		output += 'a.${name}('
		for j, _ in g.b_inps[i] {
			output += letters[i] + '_in'
			if j != g.b_inps[i].len - 1 {
				output += ', '
			}
		}
		output += ')\n'
		// push to the outputs
		for j, _ in g.b_outs[i] {
			l := letters[j]
			output += '\t\to.${l}_out.push(${l}_out)\n'
		}
		output += '\t}\n'
		output += '}\n\n'
	}
	return output
}
